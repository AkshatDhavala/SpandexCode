module fwd_core(
    input clk,
    input rst,
    
)